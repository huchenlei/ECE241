module move_validator (
  input 
  );

endmodule // move_validator
