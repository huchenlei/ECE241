module datapath (
  input
  );

endmodule // datapath
