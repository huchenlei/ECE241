module validator_b_pawn (
  input clk,
  output reg b_pawn_complete,
  input reset,
  input [2:0] piece_x, piece_y,
  input [3:0] piece_read,

  output reg [5:0] address_validator,
  output reg b_pawn_valid
  );

  // to be done later

endmodule // validator_b_pawn
