module datapath (
  input clk,
  input reset,
  input [2:0] piece_x, piece_y, // mark the selected piece
  input [2:0] box_x, box_y, // draw the select box
  input [3:0] piece_to_move
  );

endmodule // datapath
