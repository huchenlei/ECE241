module hex(hexout,   input [3:0] x;
  output [6:0]hexout;

	assign hexout[0] = (~x[3]&~x[2]&~x[1]&x[0])|(~x[3]&x[2]&~x[1]&~x[0])|(x[3]&~x[2]&x[1]&x[0])|(x[3]&x[2]&~x[1]&x[0]);
	assign hexout[1] = (~x[3]&x[2]&~x[1]&x[0])|(~x[3]&x[2]&x[1]&~x[0])|(x[3]&~x[2]&x[1]&x[0])|(x[3]&x[2]&~x[1]&~x[0])|(x[3]&x[2]&x[1]&~x[0])|(x[3]&x[2]&x[1]&x[0]);
	assign hexout[2] = (~x[3]&~x[2]&x[1]&~x[0])|(x[3]&x[2]&~x[1]&~x[0])|(x[3]&x[2]&x[1]&~x[0])|(x[3]&x[2]&x[1]&x[0]);
	assign hexout[3] = (~x[3]&~x[2]&~x[1]&x[0])|(~x[3]&x[2]&~x[1]&~x[0])|(~x[3]&x[2]&x[1]&x[0])|(x[3]&~x[2]&~x[1]&x[0])|(x[3]&~x[2]&x[1]&~x[0])|(x[3]&x[2]&x[1]&x[0]);
	assign hexout[4] = (~x[3]&~x[2]&~x[1]&x[0])|(~x[3]&~x[2]&x[1]&x[0])|(~x[3]&x[2]&~x[1]&~x[0])|(~x[3]&x[2]&~x[1]&x[0])|(~x[3]&x[2]&x[1]&x[0])|(x[3]&~x[2]&~x[1]&x[0]);
	assign hexout[5] = (~x[3]&~x[2]&~x[1]&x[0])|(~x[3]&~x[2]&x[1]&~x[0])|(~x[3]&~x[2]&x[1]&x[0])|(~x[3]&x[2]&x[1]&x[0])|(x[3]&x[2]&~x[1]&x[0]);
	assign hexout[6] = (~x[3]&~x[2]&~x[1]&~x[0])|(~x[3]&~x[2]&~x[1]&x[0])|(~x[3]&x[2]&x[1]&x[0])|(x[3]&x[2]&~x[1]&~x[0]);


endmodule
